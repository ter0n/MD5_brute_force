module brute_force_MD5(
	input logic  [31:0] MD5_A,
	input logic  [31:0] MD5_B,
	input logic  [31:0] MD5_C,
	input logic  [31:0] MD5_D,
	output logic [511:0] string_for_MD5,
	output logic 			string_ready,
	output logic [5:0]   string_length
	);

	
endmodule